module types

// This file defines the types submodule for typechecker.
