module erlang

// This file defines the erlang submodule for code generation.
