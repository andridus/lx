module generate

// This file defines the generate module.
