module erlang

// This file defines the erlang submodule for code generation.
// It includes all the files needed for Erlang code generation:
// - generator.v: Main Erlang code generator
// - expressions.v: Expression generation
// - statements.v: Statement generation
// - patterns.v: Pattern matching generation
// - formatting.v: Code formatting utilities
// - app.v: Application file generation
