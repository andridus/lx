module ast

pub struct Node {
pub:
	id       int
	kind     NodeKind
	value    string
	children []Node
	position Position
}

pub enum NodeKind {
	// Literals
	integer
	float
	string
	boolean
	atom
	nil

	// Variables
	variable_binding // x = value
	variable_ref     // x (usage)

	// Blocks
	block // do ... end or -> ... end (multiple expressions)

	// Function structure
	function
	function_body

	// Module structure
	module

	// Binary operators
	function_caller // +(a, b), *(a, b), >(a, b), etc.
	parentheses     // (expression)
}

pub struct Position {
pub:
	line   int
	column int
	file   string
}

pub struct Type {
pub:
	name   string
	params []Type
}

// Helper methods for Node
pub fn (n Node) str() string {
	return match n.kind {
		.integer { 'Int(${n.value})' }
		.float { 'Float(${n.value})' }
		.string { 'String("${n.value}")' }
		.boolean { 'Bool(${n.value})' }
		.atom { 'Atom(${n.value})' }
		.nil { 'Nil' }
		.variable_binding { 'VarBinding(${n.value})' }
		.variable_ref { 'VarRef(${n.value})' }
		.block { 'Block(${n.children.len} exprs)' }
		.function { 'Function(${n.value})' }
		.function_body { 'FunctionBody' }
		.module { 'Module' }
		.function_caller { 'FunctionCall(${n.value})' }
		.parentheses { 'Parentheses' }
	}
}

pub fn (p Position) str() string {
	return '${p.file}:${p.line}:${p.column}'
}

pub fn (t Type) str() string {
	if t.params.len == 0 {
		return t.name
	}
	params_str := t.params.map(it.str()).join(', ')
	return '${t.name}(${params_str})'
}
