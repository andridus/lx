module context

// This file defines the context submodule for code generation.
