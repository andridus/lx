module main

import parser
import lexer
import ast

// ... existing code ...
