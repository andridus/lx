module typechecker

// This file defines the typechecker module and its submodules.
