module ast

pub struct Node {
pub:
	id       int
	kind     NodeKind
	value    string
	children []Node
	position Position
}

pub enum NodeKind {
	// Literals
	integer
	float
	string
	boolean
	atom
	nil

	// Variables
	variable_binding // x = value
	variable_ref     // x (usage)
	identifier       // Generic identifier (including function args)

	// Blocks
	block // do ... end or -> ... end (multiple expressions)

	// Function structure
	function           // def function_name(args) do body end or (args) -> body
	function_parameter // function parameter definition
	lambda_expression  // fn(x) -> body end

	// Module structure
	module

	// Binary operators
	function_caller // +(a, b), *(a, b), >(a, b), etc.
	parentheses     // (expression)
	directive_call  // $print(a), $type(a)

	// List Operations
	list_literal // [1, 2, 3] ou []
	list_cons    // [head | tail]

	// Tuple Operations
	tuple_literal // {1, 2, 3} ou {}

	// Map Operations
	map_literal // %{key: value} ou %{}
	map_access  // map[key]

	// Record Operations
	record_definition // record Person { name :: string, age :: integer }
	record_field      // name :: string or name = value :: type or name = value
	record_literal    // Person{name: "João", age: 30}
	record_access     // user.name
	record_update     // %{record | campo: valor}

	// Pattern Matching
	case_expression // case expr do ... end
	case_clause     // pattern -> expression
	pattern_match   // pattern in case clause
	pattern_binding // [head | tail] = list

	// Type System
	type_alias      // type Name = Type
	type_annotation // :: Type
}

pub struct Position {
pub:
	line   int
	column int
	file   string
}

pub struct Type {
pub:
	name   string
	params []Type
}

// Helper methods for Node
pub fn (n Node) str() string {
	return '{${n.kind}, [id: ${n.id}, pos: ${n.position}], ${n.value}, ${n.children}}'
}

pub fn (p Position) str() string {
	return '${p.file}:${p.line}:${p.column}'
}

pub fn (t Type) str() string {
	if t.params.len == 0 {
		return t.name
	}
	params_str := t.params.map(it.str()).join(', ')
	return '${t.name}(${params_str})'
}

pub fn (n Node) tree_str(indent int) string {
	pad := '  '.repeat(indent)
	mut result := '${pad}{${n.kind}, [], ${n.value}, ['

	if n.children.len > 0 {
		result += '\n'
		for i, child in n.children {
			result += child.tree_str(indent + 1)
			if i < n.children.len - 1 {
				result += ','
			}
			result += '\n'
		}
		result += '${pad}]'
	} else {
		result += ']'
	}

	result += '}'
	return result
}
